`timescale 1ns / 10ps
module tb_displays_controller();




endmodule
