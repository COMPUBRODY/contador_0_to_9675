module tb_clock_divider();

endmodule
