module tb_counters_controller();

endmodule
